module imemory(reset, A, RD);

    input reset;
    input[31:0] A;
    output[31:0] RD; 

    reg[31:0] mem [1023:0];

    assign RD = (reset == 1'b0) ? {32{1'b0}} : mem[A[31:2]]; 

    
  initial begin
    $readmemh("memfile.hex",mem);
  end     



endmodule